`timescale 1ns / 1ps

module simulate_for_totaltime;

   
endmodule
