`timescale 1ns / 1ps

module turn_on_and_off(
    input clk,
    input rst,
    input power_button,  // ���ػ�����
    input left_button,
    input right_button,
    input [15:0]COUNTDOWN_TIME,
    output reg power_status, // ���ػ�״̬ (1: ����, 0: �ػ�)
    output [7:0] selection,
    output [7:0] left_time,
    output [7:0] right_time
);
    parameter LONG_PRESS_TIME = 300_000_000; // ���� 3 �� (���� 100 MHz ʱ��)
    parameter DEBOUNCE_TIME = 20_000_000;    // ȥ����ʱ 200 ms

    // �ڲ��ź�
    wire button_stable;     // ȥ����İ����ź�
    wire left_stable;       // ȥ���������ź�
    wire right_stable;      // ȥ������Ҽ��ź�
    reg [31:0] counter;     // ����������
    reg [31:0] countdown;   // ����ʱ������
    reg countdown_active;   // ����ʱ�����־
    reg is_long_press;      // ������־
    reg button_prev;        // ��һ�ΰ���״̬
    reg left_prev, right_prev;
    reg [31:0] countdown_for_time;
    // ȥ��ģ��
    debouncer #(.DEBOUNCE_TIME(DEBOUNCE_TIME)) db_power (
        .clk(clk),
        .rst(rst),
        .button_in(power_button),
        .button_out(button_stable)
    );

    debouncer #(.DEBOUNCE_TIME(DEBOUNCE_TIME)) db_left (
        .clk(clk),
        .rst(rst),
        .button_in(left_button),
        .button_out(left_stable)
    );

    debouncer #(.DEBOUNCE_TIME(DEBOUNCE_TIME)) db_right (
        .clk(clk),
        .rst(rst),
        .button_in(right_button),
        .button_out(right_stable)
    );

    // ���߼�
    always @(posedge clk or negedge rst) begin
       countdown_for_time = COUNTDOWN_TIME * 1000_0000_0;
        if (!rst) begin
            power_status <= 0; // ��ʼ״̬Ϊ�ػ�
            counter <= 0;
            is_long_press <= 0;
            countdown <= 0;
            countdown_active <= 0;
            button_prev <= 0;
            left_prev <= 0;
            right_prev <= 0;
        end else begin
            // �̰�/�����߼�
            if (button_stable) begin
                if (counter < LONG_PRESS_TIME) begin
                    counter <= counter + 1; // ��������
                end else begin
                    is_long_press <= 1; // ���Ϊ����
                end
            end else begin
                if (button_prev && !is_long_press) begin
                    power_status <= 1'b1; // �̰�����
                end else if (is_long_press) begin
                    power_status <= 1'b0; // �����ػ�
                end
                counter <= 0;
                is_long_press <= 0;
            end

            // �����߼�
            if (!power_status) begin // �ػ�״̬
                if (left_stable && !left_prev) begin
                    countdown_active <= 1;
                    countdown <= 0;
                end
                if (countdown_active && right_stable && !right_prev) begin
                    power_status <= 1; // ��� + �Ҽ� ����
                    countdown_active <= 0;
                    countdown <= 0;
                end
            end else begin // ����״̬
                if (right_stable && !right_prev) begin
                    countdown_active <= 1;
                    countdown <= 0;
                end
                if (countdown_active && left_stable && !left_prev) begin
                    power_status <= 0; // �Ҽ� + ��� �ػ�
                    countdown_active <= 0;
                    countdown <= 0;
                end
            end

            // ����ʱ�߼�
            if (countdown_active) begin
                if (countdown < countdown_for_time) begin
                    countdown <= countdown + 1;
                end else begin
                    countdown_active <= 0; // ����ʱ����
                    countdown <= 0;
                end
            end

            // ���°���״̬
            button_prev <= button_stable;
            left_prev <= left_stable;
            right_prev <= right_stable;
        end
    end
    
endmodule

// ȥ��ģ��
module debouncer #(
    parameter DEBOUNCE_TIME = 20_000_000 // ȥ����ʱ (Ĭ�� 200 ms)
)(
    input clk,
    input rst,
    input button_in,
    output reg button_out
);
    reg [24:0] counter;  // ȥ��������
    reg button_sync;     // ͬ����İ����ź�

    always @(posedge clk or negedge rst) begin
        if (!rst) begin
            counter <= 0;
            button_sync <= 0;
            button_out <= 0;
        end else begin
            button_sync <= button_in;
            if (button_sync == button_out) begin
                counter <= 0;
            end else begin
                counter <= counter + 1; // �൱�� button_sync ���źŹ���һ���ٶ���
                if (counter >= DEBOUNCE_TIME) begin
                    button_out <= button_sync;
                    counter <= 0;
                end
            end
        end
    end
endmodule
